`timescale 1 ps / 1 ps

module expr_tb ();

reg		clk;
reg		reset;
reg	[31:0]	x;
wire	[31:0]	result;

expr ex (
	.clk(clk),
	.reset(reset),
	.x(x),
	.result(result)
);

always #100 clk = ~clk;

initial
begin
	$display($time, " << Starting Simulation >> ");
	clk = 0;
	reset = 0;
	x = 32'h3f000000;
	#20000;
	$display($time, " << Simulation Complete>> ");
	$display($time, " << Simulation Complete>> ");

	$stop;
end

endmodule